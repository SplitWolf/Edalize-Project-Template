module and_gate (a,b,c);
    input a,b;
    output c;
    and (c, a, b);    
endmodule